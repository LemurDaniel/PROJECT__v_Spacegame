
module main

import gx

const (
	window_title          = 'V Spaceship Game'
	default_window_width  = 544
	default_window_height = 560
	default_background    = gx.rgb(255, 255, 255)
)